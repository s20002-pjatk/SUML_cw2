�csklearn.linear_model._logistic
LogisticRegression
q )�q}q(X   penaltyqX   l2qX   dualq�X   tolqG?6��C-X   CqG?�      X   fit_interceptq�X   intercept_scalingq	KX   class_weightq
NX   random_stateqNX   solverqX   lbfgsqX   max_iterqKdX   multi_classqX   autoqX   verboseqK X
   warm_startq�X   n_jobsqNX   l1_ratioqNX   feature_names_in_qcnumpy.core.multiarray
_reconstruct
qcnumpy
ndarray
qK �qCbq�qRq(KK�qcnumpy
dtype
qX   O8q���qRq (KX   |q!NNNJ����J����K?tq"b�]q#(X   objawyq$X   wiekq%X   chorobyq&X   wzrostq'etq(bX   n_features_in_q)KX   classes_q*hhK �q+h�q,Rq-(KK�q.hX   i8q/���q0Rq1(KX   <q2NNNJ����J����K tq3b�C               q4tq5bX   n_iter_q6hhK �q7h�q8Rq9(KK�q:hX   i4q;���q<Rq=(Kh2NNNJ����J����K tq>b�C3   q?tq@bX   coef_qAhhK �qBh�qCRqD(KKK�qEhX   f8qF���qGRqH(Kh2NNNJ����J����K tqIb�C �F��@۽|�E�}?n�>���?�A^�����qJtqKbX
   intercept_qLhhK �qMh�qNRqO(KK�qPhH�C��Z��qQtqRbX   _sklearn_versionqSX   1.0.1qTub.
��S      �sklearn.linear_model._logistic��LogisticRegression���)��}�(�penalty��l2��dual���tol�G?6��C-�C�G?�      �fit_intercept���intercept_scaling�K�class_weight�N�random_state�N�solver��lbfgs��max_iter�Kd�multi_class��auto��verbose�K �
warm_start���n_jobs�N�l1_ratio�N�feature_names_in_��numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK��h�dtype����O8�����R�(K�|�NNNJ����J����K?t�b�]�(�objawy��wiek��choroby��wzrost�et�b�n_features_in_�K�classes_�hhK ��h��R�(KK��h$�i8�����R�(K�<�NNNJ����J����K t�b�C               �t�b�n_iter_�hhK ��h��R�(KK��h$�i4�����R�(Kh9NNNJ����J����K t�b�C3   �t�b�coef_�hhK ��h��R�(KKK��h$�f8�����R�(Kh9NNNJ����J����K t�b�C �F��@۽|�E�}?n�>���?�A^������t�b�
intercept_�hhK ��h��R�(KK��hO�C��Z���t�b�_sklearn_version��1.0.1�ub.